`timescale 1ns / 1ps



module light_control1(out1,in1);

input in1;//if there is a person in the room input = 1
output out1;//if out1 is 1 turn on the light
assign out1=in1;

endmodule
