`timescale 1ns / 1ps



module water_leak_control_system(out1,in1);

input in1;//controls moisture in the basement
output out1;//if there is moisture turn of valve

assign out1=in1;

endmodule
